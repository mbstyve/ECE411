--
-- VHDL Architecture ece411.Fuck.untitled
--
-- Created:
--          by - freed2.ews (linux-a3.ews.illinois.edu)
--          at - 14:32:07 02/02/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Fuck IS
   PORT( 
      clk : IN     std_logic
   );

-- Declarations

END Fuck ;

--
ARCHITECTURE untitled OF Fuck IS
BEGIN
END ARCHITECTURE untitled;

