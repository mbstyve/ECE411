--
-- VHDL Architecture ece411.longdelay.untitled
--
-- Created:
--          by - freed2.ews (gelib-057-15.ews.illinois.edu)
--          at - 03:14:07 04/04/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY longdelay IS
   PORT( 
      F     : IN     std_logic;
      write : OUT     std_logic
   );

-- Declarations

END longdelay ;

--
ARCHITECTURE untitled OF longdelay IS
BEGIN
  write <= F after 18ns;
END ARCHITECTURE untitled;

