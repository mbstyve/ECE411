--
-- VHDL Architecture ece411.LowSig.untitled
--
-- Created:
--          by - styve1.ews (gelib-057-26.ews.illinois.edu)
--          at - 20:12:28 03/20/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;
LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY LowSig IS
   PORT( 
      A : OUT    STD_LOGIC
   );

-- Declarations

END LowSig ;

--
ARCHITECTURE untitled OF LowSig IS
BEGIN
  a <= '0';
END ARCHITECTURE untitled;

