--
-- VHDL Architecture ece411.Memory.untitled
--
-- Created:
--          by - freed2.ews (linux-a3.ews.illinois.edu)
--          at - 14:42:17 02/02/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Memory IS
   PORT( 
      ADDRESS   : IN     LC3b_word;
      DATAOUT   : IN     LC3b_word;
      MREAD_L   : IN     std_logic;
      MWRITEH_L : IN     std_logic;
      MWRITEL_L : IN     std_logic;
      RESET_L   : IN     std_logic;
      clk       : IN     std_logic;
      DATAIN    : OUT    LC3b_word;
      MRESP_H   : OUT    std_logic
   );

-- Declarations

END Memory ;

--
-- VHDL Architecture ece411.Memory.struct
--
-- Created:
--          by - freed2.ews (evrt-252-09.ews.illinois.edu)
--          at - 20:35:06 03/02/14
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;


ARCHITECTURE struct OF Memory IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL MemReadCall : std_logic;
   SIGNAL PMRESP_H    : std_logic;
   SIGNAL c_write     : std_logic;
   SIGNAL cresp_out   : std_logic;
   SIGNAL cwaitout    : std_logic;
   SIGNAL ddata       : std_logic;
   SIGNAL hitmissout  : std_logic;
   SIGNAL justdoit    : std_logic;
   SIGNAL needWB_H    : std_logic;
   SIGNAL pmaddress   : LC3B_WORD;
   SIGNAL pmdatain    : LC3B_OWORD;
   SIGNAL pmdataout   : LC3B_OWORD;
   SIGNAL pmread_l    : std_logic;
   SIGNAL pmreadstate : std_logic;
   SIGNAL pmwrite_l   : std_logic;
   SIGNAL write       : std_logic;
   SIGNAL writeback   : std_logic;


   -- Component Declarations
   COMPONENT Cache_Controller
   PORT (
      MemReadCall : IN     std_logic ;
      PMRESP_H    : IN     std_logic ;
      RESET_L     : IN     std_logic ;
      clk         : IN     std_logic ;
      hitmissout  : IN     std_logic ;
      justdoit    : IN     std_logic ;
      needWB_H    : IN     std_logic ;
      write       : IN     std_logic ;
      c_write     : OUT    std_logic ;
      cresp_out   : OUT    std_logic ;
      cwaitout    : OUT    std_logic ;
      ddata       : OUT    std_logic ;
      pmread_l    : OUT    std_logic ;
      pmreadstate : OUT    std_logic ;
      pmwrite_l   : OUT    std_logic ;
      writeback   : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Cache_Datapath
   PORT (
      ADDRESS     : IN     LC3b_word ;
      DATAOUT     : IN     LC3b_word ;
      MREAD_L     : IN     std_logic ;
      MWRITEH_L   : IN     std_logic ;
      MWRITEL_L   : IN     std_logic ;
      PMRESP_H    : IN     std_logic ;
      RESET_L     : IN     std_logic ;
      c_write     : IN     std_logic ;
      clk         : IN     std_logic ;
      cresp_out   : IN     std_logic ;
      cwaitout    : IN     std_logic ;
      ddata       : IN     std_logic ;
      pmdatain    : IN     LC3B_OWORD ;
      pmreadstate : IN     std_logic ;
      writeback   : IN     std_logic ;
      DATAIN      : OUT    LC3b_word ;
      MRESP_H     : OUT    std_logic ;
      MemReadCall : OUT    std_logic ;
      hitmissout  : OUT    std_logic ;
      needWB_H    : OUT    std_logic ;
      pmaddress   : OUT    LC3B_WORD ;
      pmdataout   : OUT    LC3B_OWORD ;
      write       : OUT    std_logic 
   );
   END COMPONENT;
   COMPONENT Physical_Memory
   PORT (
      RESET_L   : IN     std_logic ;
      clk       : IN     std_logic ;
      pmaddress : IN     LC3B_WORD ;
      pmdataout : IN     LC3B_OWORD ;
      pmread_l  : IN     std_logic ;
      pmwrite_l : IN     std_logic ;
      PMRESP_H  : OUT    std_logic ;
      pmdatain  : OUT    LC3B_OWORD 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : Cache_Controller USE ENTITY ece411.Cache_Controller;
   FOR ALL : Cache_Datapath USE ENTITY ece411.Cache_Datapath;
   FOR ALL : Physical_Memory USE ENTITY ece411.Physical_Memory;
   -- pragma synthesis_on


BEGIN

   -- Instance port mappings.
   Cache_Cont : Cache_Controller
      PORT MAP (
         MemReadCall => MemReadCall,
         PMRESP_H    => PMRESP_H,
         RESET_L     => RESET_L,
         clk         => clk,
         hitmissout  => hitmissout,
         justdoit    => justdoit,
         needWB_H    => needWB_H,
         write       => write,
         c_write     => c_write,
         cresp_out   => cresp_out,
         cwaitout    => cwaitout,
         ddata       => ddata,
         pmread_l    => pmread_l,
         pmreadstate => pmreadstate,
         pmwrite_l   => pmwrite_l,
         writeback   => writeback
      );
   Cache_DP : Cache_Datapath
      PORT MAP (
         ADDRESS     => ADDRESS,
         DATAOUT     => DATAOUT,
         MREAD_L     => MREAD_L,
         MWRITEH_L   => MWRITEH_L,
         MWRITEL_L   => MWRITEL_L,
         PMRESP_H    => PMRESP_H,
         RESET_L     => RESET_L,
         c_write     => c_write,
         clk         => clk,
         cresp_out   => cresp_out,
         cwaitout    => cwaitout,
         ddata       => ddata,
         pmdatain    => pmdatain,
         pmreadstate => pmreadstate,
         writeback   => writeback,
         DATAIN      => DATAIN,
         MRESP_H     => MRESP_H,
         MemReadCall => MemReadCall,
         hitmissout  => hitmissout,
         needWB_H    => needWB_H,
         pmaddress   => pmaddress,
         pmdataout   => pmdataout,
         write       => write
      );
   PDRAM : Physical_Memory
      PORT MAP (
         RESET_L   => RESET_L,
         clk       => clk,
         pmaddress => pmaddress,
         pmdataout => pmdataout,
         pmread_l  => pmread_l,
         pmwrite_l => pmwrite_l,
         PMRESP_H  => PMRESP_H,
         pmdatain  => pmdatain
      );

END struct;
