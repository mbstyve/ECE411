--
-- VHDL Architecture cachelib.ShifterUnit.untitled
--
-- Created:
--          by - freed2.ews (gelib-057-27.ews.illinois.edu)
--          at - 16:20:56 02/05/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY cachelib;
USE cachelib.LC3b_types.all;

ENTITY ShifterUnit IS
   PORT( 
      clk         : IN     std_logic;
      SHFTOP      : IN     LC3B_SHFTOP;
      SFTOUT      : OUT    LC3b_word;
      imm4        : IN     LC3B_NIBBLE;
      ADJ11Muxout : IN     LC3b_word
   );

-- Declarations

END ShifterUnit ;

--
ARCHITECTURE untitled OF ShifterUnit IS
BEGIN
  PROCESS (SHFTOP,ADJ11Muxout, imm4,SFTOUT)
    variable state : LC3b_word;
    variable count : integer;
  BEGIN
    case SHFTOP is
      when SHFT_SRL =>
        state := std_logic_vector("srl"(unsigned(ADJ11Muxout), to_integer(unsigned(imm4))));
      when SHFT_SLL =>
        state := std_logic_vector("sll"(unsigned(ADJ11Muxout), to_integer(unsigned(imm4))));
      when SHFT_SRA =>
        COUNT := to_integer(unsigned(imm4(3 downto 0)));
          if (imm4(3 downto 0) = "0000") then
            state := ADJ11Muxout; --Perform no shifting
          else
            state(15 - COUNT downto 0) := ADJ11Muxout(15 downto COUNT);
            state(15 downto (15 - COUNT + 1)) := (others => ADJ11Muxout(15));
          end if;
    when others =>
      state := (OTHERS => 'X');
    end case;
    SFTOUT <= state after delay_shifter;
  END PROCESS;
END ARCHITECTURE untitled;

