-- VHDL Entity ece411.EXECUTE.symbol
--
-- Created:
<<<<<<< HEAD
--          by - styve1.ews (gelib-057-20.ews.illinois.edu)
--          at - 19:31:48 04/16/14
=======
<<<<<<< HEAD
--          by - freed2.ews (gelib-057-11.ews.illinois.edu)
--          at - 22:24:23 04/15/14
=======
--          by - styve1.ews (gelib-057-14.ews.illinois.edu)
--          at - 00:56:26 04/16/14
>>>>>>> 7933d31b50383bb7b1c69148043ec0a4f94e5712
>>>>>>> d21ac329a047819d496e53151117cbb2c1e21a7b
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY EXECUTE IS
   PORT( 
      ADJ11        : IN     LC3B_WORD;
      ADJ4         : IN     LC3B_WORD;
      ADJ5         : IN     LC3B_WORD;
      ADJ6out      : IN     LC3B_WORD;
      ADJ9         : IN     lc3b_word;
      DEST         : IN     lc3b_reg;
      IMM5MuxSel   : IN     STD_LOGIC;
      JSR11        : IN     std_logic;
      RegAOut      : IN     LC3b_word;
      RegBOut      : IN     LC3B_WORD;
      SHFTOP       : IN     LC3B_SHFTOP;
      SRCA         : IN     lc3b_reg;
      SRCB         : IN     lc3b_reg;
      TRAP8        : IN     LC3B_WORD;
      control      : IN     CONTROL_WORD;
      iPC          : IN     lc3b_word  BUS;
      ADJ11_OUT    : OUT    LC3B_WORD;
      ADJ9_OUT     : OUT    LC3B_WORD;
      ALUResultout : OUT    LC3B_WORD;
      DEST_OUT     : OUT    lc3b_reg;
      JSR11_Out    : OUT    std_logic;
      RegBOut_OUT  : OUT    LC3b_word;
      SRCA_OUT     : OUT    lc3b_reg;
      SRCB_OUT     : OUT    lc3b_reg;
      TRAP8_OUT    : OUT    LC3B_WORD;
      control_out  : OUT    CONTROL_WORD;
      iPC_OUT      : OUT    lc3b_word
   );

-- Declarations

END EXECUTE ;

--
-- VHDL Architecture ece411.EXECUTE.struct
--
-- Created:
<<<<<<< HEAD
--          by - styve1.ews (gelib-057-20.ews.illinois.edu)
--          at - 19:31:48 04/16/14
=======
<<<<<<< HEAD
--          by - freed2.ews (gelib-057-11.ews.illinois.edu)
--          at - 22:24:23 04/15/14
=======
--          by - styve1.ews (gelib-057-14.ews.illinois.edu)
--          at - 00:56:26 04/16/14
>>>>>>> 7933d31b50383bb7b1c69148043ec0a4f94e5712
>>>>>>> d21ac329a047819d496e53151117cbb2c1e21a7b
--
-- Generated by Mentor Graphics' HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

LIBRARY mp3lib;

ARCHITECTURE struct OF EXECUTE IS

   -- Architecture declarations

   -- Internal signal declarations
   SIGNAL A          : STD_LOGIC;
   SIGNAL ALUAMuxSel : std_logic;
   SIGNAL ALUAMuxout : LC3B_WORD BUS;
   SIGNAL ALUMuxSel  : std_logic;
   SIGNAL ALUMuxout  : LC3B_WORD;
   SIGNAL ALUOP      : LC3B_ALUOP;
   SIGNAL ALUTrapSel : std_logic;
   SIGNAL ALUout     : LC3B_WORD;
   SIGNAL B          : LC3b_reg;
   SIGNAL F          : LC3B_WORD;
   SIGNAL F1         : LC3B_WORD;
   SIGNAL F2         : STD_LOGIC;
   SIGNAL IMM5Muxout : LC3B_WORD;
   SIGNAL ISBranch   : std_logic_vector(1 DOWNTO 0);
   SIGNAL SFTOUT     : LC3b_word;
   SIGNAL Shift      : std_logic;


   -- Component Declarations
   COMPONENT RegMux2
   PORT (
      a      : IN     LC3B_REG ;
      b      : IN     LC3B_REG ;
      Sel    : IN     std_logic ;
      Muxout : OUT    LC3B_REG 
   );
   END COMPONENT;
   COMPONENT SIGGEN111
   PORT (
      B : OUT    LC3b_reg 
   );
   END COMPONENT;
   COMPONENT Shifter
   PORT (
      SHFTOP  : IN     LC3B_SHFTOP ;
      SFTOUT  : OUT    LC3b_word ;
      RegAOut : IN     LC3b_word ;
      ADJ4    : IN     LC3B_WORD 
   );
   END COMPONENT;
   COMPONENT ctl_rip_execute
   PORT (
      control    : IN     CONTROL_WORD ;
      ALUOP      : OUT    LC3B_ALUOP ;
      ALUMuxSel  : OUT    std_logic ;
      ALUAMuxSel : OUT    std_logic ;
      Shift      : OUT    std_logic ;
      ALUTrapSel : OUT    std_logic ;
      ISBranch   : OUT    std_logic_vector (1 DOWNTO 0)
   );
   END COMPONENT;
   COMPONENT ALU
   PORT (
      A     : IN     LC3B_WORD ;
      ALUOP : IN     LC3B_ALUOP ;
      B     : IN     LC3B_WORD ;
      F     : OUT    LC3B_WORD 
   );
   END COMPONENT;
   COMPONENT AND2
   PORT (
      A : IN     STD_LOGIC ;
      B : IN     STD_LOGIC ;
      F : OUT    STD_LOGIC 
   );
   END COMPONENT;
   COMPONENT MUX2_16
   PORT (
      A   : IN     LC3B_WORD ;
      B   : IN     LC3B_WORD ;
      SEL : IN     STD_LOGIC ;
      F   : OUT    LC3B_WORD 
   );
   END COMPONENT;
   COMPONENT OR2
   PORT (
      A : IN     STD_LOGIC ;
      B : IN     STD_LOGIC ;
      F : OUT    STD_LOGIC 
   );
   END COMPONENT;

   -- Optional embedded configurations
   -- pragma synthesis_off
   FOR ALL : ALU USE ENTITY mp3lib.ALU;
   FOR ALL : AND2 USE ENTITY mp3lib.AND2;
   FOR ALL : MUX2_16 USE ENTITY mp3lib.MUX2_16;
   FOR ALL : OR2 USE ENTITY mp3lib.OR2;
   FOR ALL : RegMux2 USE ENTITY ece411.RegMux2;
   FOR ALL : SIGGEN111 USE ENTITY ece411.SIGGEN111;
   FOR ALL : Shifter USE ENTITY ece411.Shifter;
   FOR ALL : ctl_rip_execute USE ENTITY ece411.ctl_rip_execute;
   -- pragma synthesis_on


BEGIN
   -- Architecture concurrent statements
   -- HDL Embedded Text Block 1 eb1
   control_out <=control;
   DEST_OUT <= DEST;
   SRCA_OUT <= SRCA;
   SRCB_OUT <= SRCB;
   ADJ11_OUT <= ADJ11;
   ADJ9_OUT <= ADJ9;
   TRAP8_OUT <= TRAP8;
   iPC_OUT <= iPC;
   RegBOut_OUT <= RegBOut;                            


   -- Instance port mappings.
   R7Mux : RegMux2
      PORT MAP (
         a      => DEST,
         b      => B,
         Sel    => F2,
         Muxout => DEST_OUT
      );
   val7Gen : SIGGEN111
      PORT MAP (
         B => B
      );
   U_0 : Shifter
      PORT MAP (
         SHFTOP  => SHFTOP,
         SFTOUT  => SFTOUT,
         RegAOut => RegAOut,
         ADJ4    => ADJ4
      );
   execute_rip : ctl_rip_execute
      PORT MAP (
         control    => control,
         ALUOP      => ALUOP,
         ALUMuxSel  => ALUMuxSel,
         ALUAMuxSel => ALUAMuxSel,
         Shift      => Shift,
         ALUTrapSel => ALUTrapSel,
         ISBranch   => ISBranch
      );
   exALU : ALU
      PORT MAP (
         A     => ALUAMuxout,
         ALUOP => ALUOP,
         B     => ALUMuxout,
         F     => ALUout
      );
   U_3 : AND2
      PORT MAP (
         A => ISBranch(0),
         B => ISBranch(1),
         F => A
      );
   ALUAMux : MUX2_16
      PORT MAP (
         A   => RegAOut,
         B   => iPC,
         SEL => ALUAMuxSel,
         F   => ALUAMuxout
      );
   ALUMux : MUX2_16
      PORT MAP (
         A   => IMM5Muxout,
         B   => F,
         SEL => ALUMuxSel,
         F   => ALUMuxout
      );
   IMM5Mux : MUX2_16
      PORT MAP (
         A   => RegBOut,
         B   => ADJ5,
         SEL => IMM5MuxSel,
         F   => IMM5Muxout
      );
   LEAMux : MUX2_16
      PORT MAP (
         A   => ADJ6out,
         B   => F1,
         SEL => ALUAMuxSel,
         F   => F
      );
   PCoffMux : MUX2_16
      PORT MAP (
         A   => ADJ9,
         B   => TRAP8,
         SEL => ALUTrapSel,
         F   => F1
      );
   U_2 : MUX2_16
      PORT MAP (
         A   => ALUout,
         B   => SFTOUT,
         SEL => Shift,
         F   => ALUResultout
      );
   U_1 : OR2
      PORT MAP (
         A => A,
         B => ALUTrapSel,
         F => F2
      );

END struct;
