--
-- VHDL Architecture ece411.Way1.untitled
--
-- Created:
--          by - freed2.ews (gelib-057-22.ews.illinois.edu)
--          at - 15:48:50 02/13/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Way1 IS
-- Declarations

END Way1 ;

--
ARCHITECTURE untitled OF Way1 IS
BEGIN
END ARCHITECTURE untitled;

