--
-- VHDL Architecture ece411.LongNot.untitled
--
-- Created:
--          by - freed2.ews (gelib-057-15.ews.illinois.edu)
--          at - 02:08:37 04/04/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY LongNot IS
-- Declarations

END LongNot ;

--
ARCHITECTURE untitled OF LongNot IS
BEGIN
END ARCHITECTURE untitled;

